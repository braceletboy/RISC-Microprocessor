library ieee;
use ieee.std_logic_1164.all;

entity PipeRegD is
	port(
		clk, flush, freeze : in std_logic;
		
		pc_d_din, ir_d_din, ipc_d_din, r1_d_din, r2_d_din, ao_d_din : in std_logic_vector(15 downto 0);
		bm_d_din : in std_logic_vector(7 downto 0);
		
		pc_d_dout, ir_d_dout, ipc_d_dout, r1_d_dout, r2_d_dout, ao_d_dout : out std_logic_vector(15 downto 0);
		bm_d_dout : out std_logic_vector(7 downto 0);
		-- MM control signals in
		rf_a2_in_din, mem_addr_in_din, mem_din_in_din, r7_write_din, mem_write_din, ao_e_in_din : in std_logic;
		r7_din_in_din : in std_logic_vector(1 downto 0);
		-- WB control signals in
		rf_a3_in_din : in std_logic_vector(1 downto 0);
		rf_d3_in_din, reg_write_din : in std_logic;
		
		-- MM control signals out
		rf_a2_in_dout, mem_addr_in_dout, mem_din_in_dout, r7_write_dout, mem_write_dout, ao_e_in_dout : out std_logic;		
		r7_din_in_dout : out std_logic_vector(1 downto 0);
		-- WB control signals out
		rf_a3_in_dout : out std_logic_vector(1 downto 0);
		rf_d3_in_dout, reg_write_dout : out std_logic
	);
end PipeRegD;

architecture Behave of PipeRegD is
	
	signal pc_d : std_logic_vector(15 downto 0);
	signal ir_d : std_logic_vector(15 downto 0);
	signal ipc_d : std_logic_vector(15 downto 0);
	signal bm_d : std_logic_vector(7 downto 0);
	signal r1_d : std_logic_vector(15 downto 0);
	signal r2_d : std_logic_vector(15 downto 0);
	signal ao_d : std_logic_vector(15 downto 0);
	
	
	-- MM control signals
	signal rf_a2_in : std_logic;
	signal mem_addr_in : std_logic;
	signal mem_din_in : std_logic;
	signal r7_din_in : std_logic_vector(1 downto 0);
	signal r7_write : std_logic;
	signal mem_write : std_logic;
	signal ao_e_in : std_logic;
	
	-- WB control signals
	signal rf_a3_in : std_logic_vector(1 downto 0);
	signal rf_d3_in : std_logic;
	signal reg_write : std_logic;
	
begin

	process(clk, flush, freeze)
	begin
		
		if clk'event and clk = '1' then
			if flush = '1' then
				
				pc_d <= (others => '0');
				ir_d <= (others => '1');
				ipc_d <= (others => '0');
				bm_d <= (others => '0');
				r1_d <= (others => '0');
				r2_d <= (others => '0');
				ao_d <= (others => '0');
				
				
				-- MM
				rf_a2_in <= '0';
				mem_addr_in <= '0';
				mem_din_in <= '0';
				r7_din_in <= "00";
				r7_write <= '0';
				mem_write <= '0';
				ao_e_in <= '0';
				
				--WB
				rf_a3_in <= "00";
				rf_d3_in <= '0';
				reg_write <= '0';
				
			elsif freeze = '0' then
			
				pc_d <= pc_d_din;
				ir_d <= ir_d_din;
				ipc_d <= ipc_d_din;
				bm_d <= bm_d_din;
				r1_d <= r1_d_din;
				r2_d <= r2_d_din;
				ao_d <= ao_d_din;
				
				
				-- MM
				rf_a2_in <= rf_a2_in_din;
				mem_addr_in <= mem_addr_in_din;
				mem_din_in <= mem_din_in_din;
				r7_din_in <= r7_din_in_din;
				r7_write <= r7_write_din;
				mem_write <= mem_write_din;
				ao_e_in <= ao_e_in_din;
				
				-- WB
				rf_a3_in <= rf_a3_in_din;
				rf_d3_in <= rf_d3_in_din;
				reg_write <= reg_write_din;
			
			end if;
		end if;
			
		
	end process;
	
	pc_d_dout <= pc_d;
	ir_d_dout <= ir_d;
	ipc_d_dout <= ipc_d;
	bm_d_dout <= bm_d;
	r1_d_dout <= r1_d;
	r2_d_dout <= r2_d;
	ao_d_dout <= ao_d;
	
	
	-- MM
	rf_a2_in_dout <= rf_a2_in;
	mem_addr_in_dout <= mem_addr_in;
	mem_din_in_dout <= mem_din_in;
	r7_din_in_dout <= r7_din_in;
	r7_write_dout <= r7_write;
	mem_write_dout <= mem_write;
	ao_e_in_dout <= ao_e_in;
	
	-- WB
	rf_a3_in_dout <= rf_a3_in;
	rf_d3_in_dout <= rf_d3_in;
	reg_write_dout <= reg_write;

end Behave;